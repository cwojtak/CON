sal asdf false