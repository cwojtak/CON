sal asdf 256